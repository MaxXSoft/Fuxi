// a Verilog wrapper module of Fuxi
module FuxiWrapper(
  input         clk,
  input         rst,
  // interrupt requests
  input         irq_timer,
  input         irq_soft,
  input         irq_extern,
  // debug signals
  output        debug_wen,
  output [4:0]  debug_waddr,
  output [31:0] debug_wdata,
  output [31:0] debug_pc,
  // instruction AXI4 interface
  input         inst_arready,
  output        inst_arvalid,
  output [31:0] inst_araddr,
  output [3:0]  inst_arid,
  output [2:0]  inst_arsize,
  output [7:0]  inst_arlen,
  output [1:0]  inst_arburst,
  output        inst_arlock,
  output [3:0]  inst_arcache,
  output [2:0]  inst_arprot,
  output        inst_rready,
  input         inst_rvalid,
  input  [31:0] inst_rdata,
  input  [3:0]  inst_rid,
  input         inst_rlast,
  input  [1:0]  inst_rresp,
  input         inst_awready,
  output        inst_awvalid,
  output [31:0] inst_awaddr,
  output [3:0]  inst_awid,
  output [2:0]  inst_awsize,
  output [7:0]  inst_awlen,
  output [1:0]  inst_awburst,
  output        inst_awlock,
  output [3:0]  inst_awcache,
  output [2:0]  inst_awprot,
  input         inst_wready,
  output        inst_wvalid,
  output [31:0] inst_wdata,
  output [3:0]  inst_wid,
  output        inst_wlast,
  output [3:0]  inst_wstrb,
  output        inst_bready,
  input         inst_bvalid,
  input  [3:0]  inst_bid,
  input  [1:0]  inst_bresp,
  // data AXI4 interface
  input         data_arready,
  output        data_arvalid,
  output [31:0] data_araddr,
  output [3:0]  data_arid,
  output [2:0]  data_arsize,
  output [7:0]  data_arlen,
  output [1:0]  data_arburst,
  output        data_arlock,
  output [3:0]  data_arcache,
  output [2:0]  data_arprot,
  output        data_rready,
  input         data_rvalid,
  input  [31:0] data_rdata,
  input  [3:0]  data_rid,
  input         data_rlast,
  input  [1:0]  data_rresp,
  input         data_awready,
  output        data_awvalid,
  output [31:0] data_awaddr,
  output [3:0]  data_awid,
  output [2:0]  data_awsize,
  output [7:0]  data_awlen,
  output [1:0]  data_awburst,
  output        data_awlock,
  output [3:0]  data_awcache,
  output [2:0]  data_awprot,
  input         data_wready,
  output        data_wvalid,
  output [31:0] data_wdata,
  output [3:0]  data_wid,
  output        data_wlast,
  output [3:0]  data_wstrb,
  output        data_bready,
  input         data_bvalid,
  input  [3:0]  data_bid,
  input  [1:0]  data_bresp,
  // uncached AXI4 interface
  input         uncached_arready,
  output        uncached_arvalid,
  output [31:0] uncached_araddr,
  output [3:0]  uncached_arid,
  output [2:0]  uncached_arsize,
  output [7:0]  uncached_arlen,
  output [1:0]  uncached_arburst,
  output        uncached_arlock,
  output [3:0]  uncached_arcache,
  output [2:0]  uncached_arprot,
  output        uncached_rready,
  input         uncached_rvalid,
  input  [31:0] uncached_rdata,
  input  [3:0]  uncached_rid,
  input         uncached_rlast,
  input  [1:0]  uncached_rresp,
  input         uncached_awready,
  output        uncached_awvalid,
  output [31:0] uncached_awaddr,
  output [3:0]  uncached_awid,
  output [2:0]  uncached_awsize,
  output [7:0]  uncached_awlen,
  output [1:0]  uncached_awburst,
  output        uncached_awlock,
  output [3:0]  uncached_awcache,
  output [2:0]  uncached_awprot,
  input         uncached_wready,
  output        uncached_wvalid,
  output [31:0] uncached_wdata,
  output [3:0]  uncached_wid,
  output        uncached_wlast,
  output [3:0]  uncached_wstrb,
  output        uncached_bready,
  input         uncached_bvalid,
  input  [3:0]  uncached_bid,
  input  [1:0]  uncached_bresp
);

  Fuxi fuxi(
    .clock                            (clk),
    .reset                            (rst),
    // interrupt requests
    .io_irq_timer                     (irq_timer),
    .io_irq_soft                      (irq_soft),
    .io_irq_extern                    (irq_extern),
    // debug signals
    .io_debug_regWen                  (debug_wen),
    .io_debug_regWaddr                (debug_waddr),
    .io_debug_regWdata                (debug_wdata),
    .io_debug_pc                      (debug_pc),
    // instruction AXI4 interface
    .io_inst_readAddr_ready           (inst_arready),
    .io_inst_readAddr_valid           (inst_arvalid),
    .io_inst_readAddr_bits_addr       (inst_araddr),
    .io_inst_readAddr_bits_id         (inst_arid),
    .io_inst_readAddr_bits_size       (inst_arsize),
    .io_inst_readAddr_bits_len        (inst_arlen),
    .io_inst_readAddr_bits_burst      (inst_arburst),
    .io_inst_readAddr_bits_lock       (inst_arlock),
    .io_inst_readAddr_bits_cache      (inst_arcache),
    .io_inst_readAddr_bits_prot       (inst_arprot),
    .io_inst_readData_ready           (inst_rready),
    .io_inst_readData_valid           (inst_rvalid),
    .io_inst_readData_bits_data       (inst_rdata),
    .io_inst_readData_bits_id         (inst_rid),
    .io_inst_readData_bits_last       (inst_rlast),
    .io_inst_readData_bits_resp       (inst_rresp),
    .io_inst_writeAddr_ready          (inst_awready),
    .io_inst_writeAddr_valid          (inst_awvalid),
    .io_inst_writeAddr_bits_addr      (inst_awaddr),
    .io_inst_writeAddr_bits_id        (inst_awid),
    .io_inst_writeAddr_bits_size      (inst_awsize),
    .io_inst_writeAddr_bits_len       (inst_awlen),
    .io_inst_writeAddr_bits_burst     (inst_awburst),
    .io_inst_writeAddr_bits_lock      (inst_awlock),
    .io_inst_writeAddr_bits_cache     (inst_awcache),
    .io_inst_writeAddr_bits_prot      (inst_awprot),
    .io_inst_writeData_ready          (inst_wready),
    .io_inst_writeData_valid          (inst_wvalid),
    .io_inst_writeData_bits_data      (inst_wdata),
    .io_inst_writeData_bits_id        (inst_wid),
    .io_inst_writeData_bits_last      (inst_wlast),
    .io_inst_writeData_bits_strb      (inst_wstrb),
    .io_inst_writeResp_ready          (inst_bready),
    .io_inst_writeResp_valid          (inst_bvalid),
    .io_inst_writeResp_bits_id        (inst_bid),
    .io_inst_writeResp_bits_resp      (inst_bresp),
    // data AXI4 interface
    .io_data_readAddr_ready           (data_arready),
    .io_data_readAddr_valid           (data_arvalid),
    .io_data_readAddr_bits_addr       (data_araddr),
    .io_data_readAddr_bits_id         (data_arid),
    .io_data_readAddr_bits_size       (data_arsize),
    .io_data_readAddr_bits_len        (data_arlen),
    .io_data_readAddr_bits_burst      (data_arburst),
    .io_data_readAddr_bits_lock       (data_arlock),
    .io_data_readAddr_bits_cache      (data_arcache),
    .io_data_readAddr_bits_prot       (data_arprot),
    .io_data_readData_ready           (data_rready),
    .io_data_readData_valid           (data_rvalid),
    .io_data_readData_bits_data       (data_rdata),
    .io_data_readData_bits_id         (data_rid),
    .io_data_readData_bits_last       (data_rlast),
    .io_data_readData_bits_resp       (data_rresp),
    .io_data_writeAddr_ready          (data_awready),
    .io_data_writeAddr_valid          (data_awvalid),
    .io_data_writeAddr_bits_addr      (data_awaddr),
    .io_data_writeAddr_bits_id        (data_awid),
    .io_data_writeAddr_bits_size      (data_awsize),
    .io_data_writeAddr_bits_len       (data_awlen),
    .io_data_writeAddr_bits_burst     (data_awburst),
    .io_data_writeAddr_bits_lock      (data_awlock),
    .io_data_writeAddr_bits_cache     (data_awcache),
    .io_data_writeAddr_bits_prot      (data_awprot),
    .io_data_writeData_ready          (data_wready),
    .io_data_writeData_valid          (data_wvalid),
    .io_data_writeData_bits_data      (data_wdata),
    .io_data_writeData_bits_id        (data_wid),
    .io_data_writeData_bits_last      (data_wlast),
    .io_data_writeData_bits_strb      (data_wstrb),
    .io_data_writeResp_ready          (data_bready),
    .io_data_writeResp_valid          (data_bvalid),
    .io_data_writeResp_bits_id        (data_bid),
    .io_data_writeResp_bits_resp      (data_bresp),
    // uncached AXI4 interface
    .io_uncached_readAddr_ready       (uncached_arready),
    .io_uncached_readAddr_valid       (uncached_arvalid),
    .io_uncached_readAddr_bits_addr   (uncached_araddr),
    .io_uncached_readAddr_bits_id     (uncached_arid),
    .io_uncached_readAddr_bits_size   (uncached_arsize),
    .io_uncached_readAddr_bits_len    (uncached_arlen),
    .io_uncached_readAddr_bits_burst  (uncached_arburst),
    .io_uncached_readAddr_bits_lock   (uncached_arlock),
    .io_uncached_readAddr_bits_cache  (uncached_arcache),
    .io_uncached_readAddr_bits_prot   (uncached_arprot),
    .io_uncached_readData_ready       (uncached_rready),
    .io_uncached_readData_valid       (uncached_rvalid),
    .io_uncached_readData_bits_data   (uncached_rdata),
    .io_uncached_readData_bits_id     (uncached_rid),
    .io_uncached_readData_bits_last   (uncached_rlast),
    .io_uncached_readData_bits_resp   (uncached_rresp),
    .io_uncached_writeAddr_ready      (uncached_awready),
    .io_uncached_writeAddr_valid      (uncached_awvalid),
    .io_uncached_writeAddr_bits_addr  (uncached_awaddr),
    .io_uncached_writeAddr_bits_id    (uncached_awid),
    .io_uncached_writeAddr_bits_size  (uncached_awsize),
    .io_uncached_writeAddr_bits_len   (uncached_awlen),
    .io_uncached_writeAddr_bits_burst (uncached_awburst),
    .io_uncached_writeAddr_bits_lock  (uncached_awlock),
    .io_uncached_writeAddr_bits_cache (uncached_awcache),
    .io_uncached_writeAddr_bits_prot  (uncached_awprot),
    .io_uncached_writeData_ready      (uncached_wready),
    .io_uncached_writeData_valid      (uncached_wvalid),
    .io_uncached_writeData_bits_data  (uncached_wdata),
    .io_uncached_writeData_bits_id    (uncached_wid),
    .io_uncached_writeData_bits_last  (uncached_wlast),
    .io_uncached_writeData_bits_strb  (uncached_wstrb),
    .io_uncached_writeResp_ready      (uncached_bready),
    .io_uncached_writeResp_valid      (uncached_bvalid),
    .io_uncached_writeResp_bits_id    (uncached_bid),
    .io_uncached_writeResp_bits_resp  (uncached_bresp)
  );

endmodule
